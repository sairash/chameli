module main


import lexer

fn main() {
	println(lexer.Lex.new(""))
}
