module lexer

import token
